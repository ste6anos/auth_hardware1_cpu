`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:30:50 01/04/2022 
// Design Name: 
// Module Name:    decoder5to32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module decoder5to32(
          input [4:0] a,
			 input en, 
			 output [31:0] decout
    );
   reg[31:0] out;
	assign decout= out;
   always @(*)
	begin
	 if(en) begin
	   case(a) 
	     0:  out = 32'b00000000000000000000000000000001;
	     1:  out = 32'b00000000000000000000000000000010;
	     2:  out = 32'b00000000000000000000000000000100;
	     3:  out = 32'b00000000000000000000000000001000;
		  4:  out = 32'b00000000000000000000000000010000;
		  5:  out = 32'b00000000000000000000000000100000;
		  6:  out = 32'b00000000000000000000000001000000;
	     7:  out = 32'b00000000000000000000000010000000;
	     8:  out = 32'b00000000000000000000000100000000;
	     9:  out = 32'b00000000000000000000001000000000;
		 10:  out = 32'b00000000000000000000010000000000;
		 11:  out = 32'b00000000000000000000100000000000;
		 12:  out = 32'b00000000000000000001000000000000;
	    13:  out = 32'b00000000000000000010000000000000;
	    14:  out = 32'b00000000000000000100000000000000;
	    15:  out = 32'b00000000000000001000000000000000;
		 16:  out = 32'b00000000000000010000000000000000;
		 17:  out = 32'b00000000000000100000000000000000;
	    18:  out = 32'b00000000000001000000000000000000;
	    19:  out = 32'b00000000000010000000000000000000;
	    20:  out = 32'b00000000000100000000000000000000;
		 21:  out = 32'b00000000001000000000000000000000;
		 22:  out = 32'b00000000010000000000000000000000;
		 23:  out = 32'b00000000100000000000000000000000;
	    24:  out = 32'b00000001000000000000000000000000;
	    25:  out = 32'b00000010000000000000000000000000;
	    26:  out = 32'b00000100000000000000000000000000;
		 27:  out = 32'b00001000000000000000000000000000;
		 28:  out = 32'b00010000000000000000000000000000;
		 29:  out = 32'b00100000000000000000000000000000;
		 30:  out = 32'b01000000000000000000000000000000;
		 31:  out = 32'b10000000000000000000000000000000;
      default out=0;
		endcase
    end
	 else 
	  out =0;
   end
	
	
	
	

endmodule
